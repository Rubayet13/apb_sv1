`include "apb_slave.svp"
`include "apb_interface.sv"
`include "apb_monitor.sv"
`include "apb_driver.sv"
`include "apb_agent.sv"
`include "apb_scb.sv"
`include "apb_env.sv"
`include "apb_test.sv"
