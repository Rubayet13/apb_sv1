class apb_scb; 
	function new (string name = "apb_scb", virtual apb_intf INTF);
		$display ("%s is created", name);
	endfunction 
endclass 
